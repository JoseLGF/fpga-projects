H���   о��   X҂�   ���   h���   ���   x ��    4��   �G��   [��   �n��    ���   ����   0���   ����   @Ѓ�   ���   P���   �
��   `��   �1��   pE��   �X��   �l��   ���   ����   ���   ����   (΄�   ���   8���   ���   H��   �/��   XC��   �V��   hj��   �}��   x���    ���   ����   ̅�   �߅�    ��   ���   0��   �-��   @A��   �T��   Ph��   �{��   `���   袆�   p���   �Ɇ�   �݆�   ��   ���   ��   �+��   (?��   �R��   8f��   �y��   H���   Р��   X���   �Ǉ�   hۇ�   ���   x��    ��   �)��   =��   �P��    d��   �w��   0���   ����   @���   �ň�   Pو�   ���   ` ��   ���   p'��   �:��   �N��   b��   �u��   ���   ����   (���   �É�   8׉�   ���   H���   ���   X%��   �8��   hL��   �_��   xs��    ���   ����   ���   ����    Պ�   ���   0���   ���   @#��   �6��   PJ��   �]��   `q��   脋�   p���   ����   ����   Ӌ�   ���   ���   ���   (!��   �4��   8H��   �[��   Ho��   Ђ��   X���   ੌ�   h���   �Ќ�   x��    ���   ���   ��   �2��    F��   �Y��   0m��   ����   @���   ȧ��   P���   �΍�   `��   ����   p	��   ���   �0��   D��   �W��   k��   �~��   (���   ����   8���   �̎�   H���   ���   X��   ���   h.��   �A��   xU��    i��   �|��   ���   ����    ���   �ʏ�   0ޏ�   ���   @��   ���   P,��   �?��   `S��   �f��   pz��   ����   ����   ���   �Ȑ�   ܐ�   ���   (��   ���   8*��   �=��   HQ��   �d��   Xx��   ����   h���   ��   xƑ�    ڑ�   ���   ��   ���    (��   �;��   0O��   �b��   @v��   ȉ��   P���   ذ��   `Ē�   �ג�   p��   ����   ���   &��   �9��   M��   �`��   (t��   ����   8���   ����   H�   �Փ�   X��   ����   h��   �#��   x7��    K��   �^��   r��   ����    ���   ����   0���   �Ӕ�   @��   ����   P��   �!��   `5��   �H��   p\��   �o��   ����   ���   ����   ���   �ѕ�   (��   ����   8��   ���   H3��   �F��   XZ��   �m��   h���   ��   x���    ���   �ϖ�   ��   ����    
��   ���   01��   �D��   @X��   �k��   P��   ؒ��   `���   蹗�   p͗�   ����   ����   ��   ���   /��   �B��   (V��   �i��   8}��   ����   H���   з��   X˘�   �ޘ�   h��   ���   x��    -��   �@��   T��   �g��    {��   ����   0���   ����   @ə�   �ܙ�   P��   ���   `��   �*��   p>��   �Q��   �e��   y��   ����   ���   ����   (ǚ�   �ښ�   8��   ���   H��   �(��   X<��   �O��   hc��   �v��   x���    ���   ����   ś�   �؛�    ��   ����   0��   �&��   @:��   �M��   Pa��   �t��   `���   蛜�   p���   ��   �֜�   ��   ����   ��   �$��   (8��   �K��   8_��   �r��   H���   Й��   X���   ����   hԝ�   ���   x���    ��   �"��   6��   �I��    ]��   �p��   0���   ����   @���   Ⱦ��   PҞ�   ���   `���   ���   p ��   �3��   �G��   [��   �n��   ���   ����   (���   ����   8П�   ���   H���   �
��   X��   �1��   hE��   �X��   xl��   